module dmac_data_mover (
	input s_axi_aclk,
	input s_axi_aresetn,

	input [C_ID_WIDTH-1:0] request_id,
	output [C_ID_WIDTH-1:0] response_id,
	input sync_id,
	input eot,

	input enable,
	output reg enabled,

	output s_axi_ready,
	input s_axi_valid,
	input [C_DATA_WIDTH-1:0] s_axi_data,

	input m_axi_ready,
	output m_axi_valid,
	output [C_DATA_WIDTH-1:0] m_axi_data,
	output m_axi_last,

	input req_valid,
	output reg req_ready,
	input [3:0] req_last_burst_length
);

parameter C_ID_WIDTH = 3;
parameter C_DATA_WIDTH = 64;
parameter C_DISABLE_WAIT_FOR_ID = 1;

`include "inc_id.v"

reg [3:0] last_burst_length;
reg [C_ID_WIDTH-1:0] id = 'h00;
reg [C_ID_WIDTH-1:0] id_next;
reg [3:0] beat_counter = 'h00;
wire [3:0] beat_counter_next;
wire last;
reg pending_burst;

assign response_id = id;

assign beat_counter_next = s_axi_ready && s_axi_valid ? beat_counter + 1'b1 : beat_counter;
assign last = beat_counter == (eot ? last_burst_length : 4'hf);

assign s_axi_ready = m_axi_ready & pending_burst & ~req_ready;
assign m_axi_valid = s_axi_valid & pending_burst & ~req_ready;
assign m_axi_data = s_axi_data;
assign m_axi_last = last;

always @(posedge s_axi_aclk) begin
	if (s_axi_aresetn == 1'b0) begin
		enabled <= 1'b0;
	end else begin
		if (enable) begin
			enabled <= 1'b1;
		end else begin
			if (C_DISABLE_WAIT_FOR_ID == 0) begin
				// We are not allowed to just deassert valid, so wait until the
				// current beat has been accepted
				if (~s_axi_valid || m_axi_ready)
					enabled <= 1'b0;
			end else begin
				// For memory mapped AXI busses we have to complete all pending
				// burst requests before we can disable the data mover.
				if (response_id == request_id)
					enabled <= 1'b0;
			end
		end
	end
end

always @(posedge s_axi_aclk) begin
	if (s_axi_aresetn == 1'b0) begin
		beat_counter <= 'h0;
		req_ready <= 1'b1;
	end else begin
		if (~enabled) begin
			req_ready <= 1'b1;
		end else if (req_ready) begin
			if (req_valid && enabled) begin
				last_burst_length <= req_last_burst_length;
				req_ready <= 1'b0;
				beat_counter <= 'h0;
			end
		end else if (s_axi_ready && s_axi_valid) begin
			if (last && eot)
				req_ready <= 1'b1;
			beat_counter <= beat_counter + 1'b1;
		end
	end
end

always @(*)
begin
	if ((s_axi_ready && s_axi_valid && last) ||
		(sync_id && id != request_id))
		id_next <= inc_id(id);
	else
		id_next <= id;
end

always @(posedge s_axi_aclk) begin
	if (s_axi_aresetn == 1'b0) begin
		id <= 'h0;
	end else begin
		id <= id_next;
		pending_burst <= id_next != request_id;
	end
end

endmodule
